function int fac_function (input int m,n);
	int fac_function = 1;
	for(int i =1; i< m+n+1; i++)
		fac_function *= i;
endfunction
